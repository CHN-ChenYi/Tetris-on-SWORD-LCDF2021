`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:    15:31:35 01/10/2021
// Design Name:
// Module Name:    Rotate
// Project Name:
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
module Rotate(
         input wire clk,
         input wire [0:15] float, // float blocks' status
         input wire direction, // 0 for clockwise
         output wire [0:15] new_float // after rotation
       );


endmodule
